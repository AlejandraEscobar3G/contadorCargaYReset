library verilog;
use verilog.vl_types.all;
entity contadorEstado_vlg_vec_tst is
end contadorEstado_vlg_vec_tst;
